`define FUNCT_ADD 6'b100000
`define FUNCT_SUB 6'b100010
`define FUNCT_AND 6'b100100
`define FUNCT_OR 6'b100101
`define FUNCT_SLT 6'b101010

`define OP_R 6'b000000
`define OP_LW 6'b100011
`define OP_SW 6'b101011
`define OP_BEQ 6'b000100
`define OP_BNE 6'b000101
`define OP_ADDI 6'b001000
`define OP_SLTI 6'b001010
`define OP_ORI 6'b001101
`define OP_ANDI 6'b001100
`define OP_J 6'b000010